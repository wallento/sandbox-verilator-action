module A;
    wire [1:0] a;

    assign a = 2'b01;
endmodule
